��/  K��@AZ�����"SƤ`��g�o[j#ƽ�n-1��͈�P�Ǜ�*e�c�1��E#nT-�}����](0��'d���a�n�ƪ��H�.�1_�`1(WB>M�{*3��J�{|�S�&|}�@~H��c�9O�t�����}�n葥����29iY�IX����V�W|D&��1�^k��}��Tl�/*֍�����NX|���?�Q���`�C���q�43k�{tn�cVo $�$��q�W$�-��re �&{�s�B��>(y/nV���O���.s� �@J��Q�(��A@�C�q�*{������4��w�JL��y:���ҕ�@w�$�\��z��,��=0#�̑���0��Z��+�
��znY�+b��]Q���"�AX��s�3L̸e؉�9j�5�)��(=@NG���a�+R�q8�'R���^	d�$!���@�Q���������V���WѤ^��hW�T&9g�>v���ۡ�B�s�O�"� e*��t�7ݴ����EU��m��u���@�(����:<�$�|�
��M��e|#ee��	VD�u��B�%>�X��w �Q��&L{/Ԍ`���HL~�<�Os��l�l^8x(�\�5e����{�� H]����?n�W��l �=�d:X�[@s��D�^̢��LΗ�o�{��_�!<L;��2���fT�<$ʏ�2�{F�jG����&�~�k��ZS�;I9��(�� ����c�C��c�!F\]4wHǘHZ������h�FJcw��XD���h˹�U+���b���ei��n�
��p1/�dcK�������y���J~_'՝[�%�md+�)�d�e�Q��suy�$�k��Id�~{�E~���@��=���,B��И�u��?�BA�J�7w�V����Z58'<�;�PIaf���&�f�-�c`�U$���p�ي�����ݥS�R���)fZf��-$�Vj0G�u�������q�g�~���M����0���$wG�I�	����I��+0�	�� ��B�_l���"|;�Ԯ�RՃ�XZ
��=C�/BC���ZU���07�zI1�9�bK#����`���8�0Kx}7��\0��D�c�����HǵI���T�)���Ѯ�����&��j�0�*vĎ�:�vR�5Q�yw]�U�x�86w.lˋ{ M��Q���ͣ�������k�w"AY7)���5l��z���ٵ^�E(�ji�I�Qȉ�ˍ��ǵ$��XU})wa�������wc,2��t﷠��P@T���q�#��ͅZ�+��9�֧!���ϣJo�m�eMUX��"�	��n���c��r|g��hӮ��XU SP�Z&�v�Sq�F�ű�Jc�w�X������K���<���ϡ�CA��
�XS�/	O�dh�oV>k��u	���xAo��a�MK��
���6��D���Zܣ�}={*� �ּ�p�i�7:Ӌ�C]����NG` 7=�ea1^"�5�wp������^h��ϋT�)�6��y��@�!���=�n���4�yGq�%��8��;�R��ru��#�����A@���ׂB�ڞN`z~Ujw%p��N<�9����/��J�.qI��A#�wh�NrSW�$�k,��Ϙ�)s�r���3�� �h�T���-�=�Z�b����E�����^ݮ�<��X�xJ.����}<�h{���ߌDC2��NN���s?�;m�0�T*j)��y��0��S) ���g>�	��ȇҟ;���RB�OU.��ŏ���Y<T��uQ:��4��i&�,�0fi�R��m(~�n�)��$�->d�M�����p����f��/M�U�o�����0�IqĶ��v�����!�����E�Q�JNS�(���	��Έ�I��9 $e�異q?H��-Oπ#��^��/Y��)xFᯊGq��l@m^%�*���,��($���;6���M��v�gb)3�w�� L�B�Z]���y��Ze>��
�I�������6U��/c��i�E�6�*���	��B
"�f���_���Eȫ������/��H���jٌR��w�*X�K#�T�߄9G}o��Ci�{2�l@Ԥ��gч�w�̔�~�H}k.����n"\�/!Z�z:�sY��=��椶�Źr���K�o�B�뗖!<��D�/Wy��/s���0�e�5P3?��f}��ʂxǍ�_�%B�+Y�*W��<��YX�Il�=X�h)n7'څ&����0S�E������O�9��.L�5Q7��og����
wyrЅ�J�Dk���W�`��7�$gT�����r�!������|���ru��l��it�ӳ�z����Ɗ��mC����6J?z]ߒ�!e��jM���q��:�1��e�?-b�@"�71��{���\Ì�<�u;�����s���:-�aJ�iL�6���H3�$��4��m֋b��[#��W���c��?��`���p���]y��bd�޼<��v���&D,�m1��6�Ou?ݯѶa�(���Z!²vv�J�fO�F��\�]�߿2[�jN���Lu�$Ni����3���� ����9:3��!O���J>�U)/�8���Li���C�E�����-H��?>!�$H�㥪}+� �r�H��{���I��A�@�. �}V�7t��T��a`x6���͋��y����,Ԁ��O�`��H��[b���"E��_����,v�k�v�ᏸ����Ʉ���T�Z���Xr��l�J��4D�̕��Cd4("oi���7<	>��6�^���뽕��pq��x�� ��K���aG���RF?m<|V���M��B2C"��w�0m�Fa<Cٖ��tT�kU������*���M��!����0��֝�Ϙ�yG���v�'�oNC�A'�����"qj��#��
І��j�o���Ax��N{s;���?	~?u�3J�b�x���+v��_�*���WQ���4�u%t$�d�������/���+]��cBx� ���c���
xHG1�����g����tU$m�i�3���!��m��3�J�����S^t�.5��MZo'/�w�/���Goi
��tz�����-��5RC"�.-[Q:�Z���K٠#SI�,�a_m��5_Q���P�*ZPQo1�<��o���r�Cf<���� a�{�u���8	����f��f"�b�@B�AS*yV�C���0�r]-���]��~q���p� �ZScd�e@h(%�'e�88Һ���S��L�H{�e�D�b� 硫x���VY�sH��)ŝ2v�VQ�����UhvÖ��>�_�é�48l���?1��X��2��C9����M���4@AHj���V�}l�F!74�<z�hN-1��;"E��G^7昌 �bT�2�� �5D?��9Ψ�t{����D��}6�;��>hA����ܣ��E���
�*c*�ק�/8�u�yd74���&����_��^�p��
�I��}S�IK|�`��UH�:4�Q�S`
����yy"�*�0��,d�V��[����Ym����Ef�58�0���0b!���������+J�ڥ𠯵O$�
,t8G\��UUʑv֡B�δ��x�?�3�g#�_������|0�hKPe�.��L��l0i��N?�X��ˠs�쵲��O�9{iͩ7��MqSvT��a��Nsgs��~#�j���G	I�_j����fja��Ġ3�5/j綃Z���4t�K0P���0����T��U��ZO8�[���I���Vy���_��Z���)�[бU*��(OJ��07�i/��G�a��l\�m:�r�C���Τe2�K����=^�Ake,8��ƹG�2�}�f��,�>-Ͱ�e`�}�ܐ`�K����y���Y�����7W�2{$����D��m���M?E����4�3��1�g��fI%�#�u�F��&:��K7}����ݮ�3_����	}:?�b�y�7@U�\0%߇H'��̪S��d�!��>w�W%��?��D��D9��U��\�����	��!KU�p-��v8�fx��n}�8�p��g4�w��|�o|"Ɨ���yE�'awm�" Z�A����Bϳ&s�ͳh��>�?��C�r-*U<����p���>�rA-�+�g7x����`	mB|��������n�j��X�Wv���'�	�L��n˼�� �ube@�X(PU>?��_�.��oXn��81�d_�F,�!A��30Iц�1J��g�FX�p�Һ�=�ʳ8��� ��N��*��!L�>c0�_+��,.{aH��C�i
��݄>ϛ��K�����d�4�J��Pq�Ĳ�j���݆�{�%��7D!�4��b�-l��ϒ��-�ڿ߻�X�2PZ&�Ie�|Tb(�0�v��:����ϻ���{�ȥ�N%Q�۬'�f�x�X���Q�n؃ݙ؟S��� �h�E!�����Ř�)�E�OT0���Ǽc��iP�m�rg�Gҹ{����^N��L;?�}����